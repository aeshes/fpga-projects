module sine_signal(
    input logic clk,
    output logic [0:7] signal
);

    logic [0:7] counter;

    sawtooth_signal sawtooth(clk, counter);

    always_ff @(posedge clk)
    begin
        case (counter)
            8'b00000000: signal <= 8'b01111111;
            8'b00000001: signal <= 8'b10000010;
            8'b00000010: signal <= 8'b10000101;
            8'b00000011: signal <= 8'b10001000;
            8'b00000100: signal <= 8'b10001011;
            8'b00000101: signal <= 8'b10001110;
            8'b00000110: signal <= 8'b10010001;
            8'b00000111: signal <= 8'b10010100;
            8'b00001000: signal <= 8'b10010111;
            8'b00001001: signal <= 8'b10011010;
            8'b00001010: signal <= 8'b10011101;
            8'b00001011: signal <= 8'b10100000;
            8'b00001100: signal <= 8'b10100011;
            8'b00001101: signal <= 8'b10100110;
            8'b00001110: signal <= 8'b10101001;
            8'b00001111: signal <= 8'b10101100;
            8'b00010000: signal <= 8'b10101111;
            8'b00010001: signal <= 8'b10110010;
            8'b00010010: signal <= 8'b10110101;
            8'b00010011: signal <= 8'b10111000;
            8'b00010100: signal <= 8'b10111010;
            8'b00010101: signal <= 8'b10111101;
            8'b00010110: signal <= 8'b11000000;
            8'b00010111: signal <= 8'b11000010;
            8'b00011000: signal <= 8'b11000101;
            8'b00011001: signal <= 8'b11001000;
            8'b00011010: signal <= 8'b11001010;
            8'b00011011: signal <= 8'b11001101;
            8'b00011100: signal <= 8'b11001111;
            8'b00011101: signal <= 8'b11010001;
            8'b00011110: signal <= 8'b11010100;
            8'b00011111: signal <= 8'b11010110;
            8'b00100000: signal <= 8'b11011000;
            8'b00100001: signal <= 8'b11011010;
            8'b00100010: signal <= 8'b11011101;
            8'b00100011: signal <= 8'b11011111;
            8'b00100100: signal <= 8'b11100001;
            8'b00100101: signal <= 8'b11100011;
            8'b00100110: signal <= 8'b11100101;
            8'b00100111: signal <= 8'b11100110;
            8'b00101000: signal <= 8'b11101000;
            8'b00101001: signal <= 8'b11101010;
            8'b00101010: signal <= 8'b11101011;
            8'b00101011: signal <= 8'b11101101;
            8'b00101100: signal <= 8'b11101111;
            8'b00101101: signal <= 8'b11110000;
            8'b00101110: signal <= 8'b11110001;
            8'b00101111: signal <= 8'b11110011;
            8'b00110000: signal <= 8'b11110100;
            8'b00110001: signal <= 8'b11110101;
            8'b00110010: signal <= 8'b11110110;
            8'b00110011: signal <= 8'b11110111;
            8'b00110100: signal <= 8'b11111000;
            8'b00110101: signal <= 8'b11111001;
            8'b00110110: signal <= 8'b11111010;
            8'b00110111: signal <= 8'b11111010;
            8'b00111000: signal <= 8'b11111011;
            8'b00111001: signal <= 8'b11111100;
            8'b00111010: signal <= 8'b11111100;
            8'b00111011: signal <= 8'b11111101;
            8'b00111100: signal <= 8'b11111101;
            8'b00111101: signal <= 8'b11111101;
            8'b00111110: signal <= 8'b11111101;
            8'b00111111: signal <= 8'b11111101;
            8'b01000000: signal <= 8'b11111110;
            8'b01000001: signal <= 8'b11111101;
            8'b01000010: signal <= 8'b11111101;
            8'b01000011: signal <= 8'b11111101;
            8'b01000100: signal <= 8'b11111101;
            8'b01000101: signal <= 8'b11111101;
            8'b01000110: signal <= 8'b11111100;
            8'b01000111: signal <= 8'b11111100;
            8'b01001000: signal <= 8'b11111011;
            8'b01001001: signal <= 8'b11111010;
            8'b01001010: signal <= 8'b11111010;
            8'b01001011: signal <= 8'b11111001;
            8'b01001100: signal <= 8'b11111000;
            8'b01001101: signal <= 8'b11110111;
            8'b01001110: signal <= 8'b11110110;
            8'b01001111: signal <= 8'b11110101;
            8'b01010000: signal <= 8'b11110100;
            8'b01010001: signal <= 8'b11110011;
            8'b01010010: signal <= 8'b11110001;
            8'b01010011: signal <= 8'b11110000;
            8'b01010100: signal <= 8'b11101111;
            8'b01010101: signal <= 8'b11101101;
            8'b01010110: signal <= 8'b11101011;
            8'b01010111: signal <= 8'b11101010;
            8'b01011000: signal <= 8'b11101000;
            8'b01011001: signal <= 8'b11100110;
            8'b01011010: signal <= 8'b11100101;
            8'b01011011: signal <= 8'b11100011;
            8'b01011100: signal <= 8'b11100001;
            8'b01011101: signal <= 8'b11011111;
            8'b01011110: signal <= 8'b11011101;
            8'b01011111: signal <= 8'b11011010;
            8'b01100000: signal <= 8'b11011000;
            8'b01100001: signal <= 8'b11010110;
            8'b01100010: signal <= 8'b11010100;
            8'b01100011: signal <= 8'b11010001;
            8'b01100100: signal <= 8'b11001111;
            8'b01100101: signal <= 8'b11001101;
            8'b01100110: signal <= 8'b11001010;
            8'b01100111: signal <= 8'b11001000;
            8'b01101000: signal <= 8'b11000101;
            8'b01101001: signal <= 8'b11000010;
            8'b01101010: signal <= 8'b11000000;
            8'b01101011: signal <= 8'b10111101;
            8'b01101100: signal <= 8'b10111010;
            8'b01101101: signal <= 8'b10111000;
            8'b01101110: signal <= 8'b10110101;
            8'b01101111: signal <= 8'b10110010;
            8'b01110000: signal <= 8'b10101111;
            8'b01110001: signal <= 8'b10101100;
            8'b01110010: signal <= 8'b10101001;
            8'b01110011: signal <= 8'b10100110;
            8'b01110100: signal <= 8'b10100011;
            8'b01110101: signal <= 8'b10100000;
            8'b01110110: signal <= 8'b10011101;
            8'b01110111: signal <= 8'b10011010;
            8'b01111000: signal <= 8'b10010111;
            8'b01111001: signal <= 8'b10010100;
            8'b01111010: signal <= 8'b10010001;
            8'b01111011: signal <= 8'b10001110;
            8'b01111100: signal <= 8'b10001011;
            8'b01111101: signal <= 8'b10001000;
            8'b01111110: signal <= 8'b10000101;
            8'b01111111: signal <= 8'b10000010;
            8'b10000000: signal <= 8'b01111111;
            8'b10000001: signal <= 8'b01111011;
            8'b10000010: signal <= 8'b01111000;
            8'b10000011: signal <= 8'b01110101;
            8'b10000100: signal <= 8'b01110010;
            8'b10000101: signal <= 8'b01101111;
            8'b10000110: signal <= 8'b01101100;
            8'b10000111: signal <= 8'b01101001;
            8'b10001000: signal <= 8'b01100110;
            8'b10001001: signal <= 8'b01100011;
            8'b10001010: signal <= 8'b01100000;
            8'b10001011: signal <= 8'b01011101;
            8'b10001100: signal <= 8'b01011010;
            8'b10001101: signal <= 8'b01010111;
            8'b10001110: signal <= 8'b01010100;
            8'b10001111: signal <= 8'b01010001;
            8'b10010000: signal <= 8'b01001110;
            8'b10010001: signal <= 8'b01001011;
            8'b10010010: signal <= 8'b01001000;
            8'b10010011: signal <= 8'b01000101;
            8'b10010100: signal <= 8'b01000011;
            8'b10010101: signal <= 8'b01000000;
            8'b10010110: signal <= 8'b00111101;
            8'b10010111: signal <= 8'b00111011;
            8'b10011000: signal <= 8'b00111000;
            8'b10011001: signal <= 8'b00110101;
            8'b10011010: signal <= 8'b00110011;
            8'b10011011: signal <= 8'b00110000;
            8'b10011100: signal <= 8'b00101110;
            8'b10011101: signal <= 8'b00101100;
            8'b10011110: signal <= 8'b00101001;
            8'b10011111: signal <= 8'b00100111;
            8'b10100000: signal <= 8'b00100101;
            8'b10100001: signal <= 8'b00100011;
            8'b10100010: signal <= 8'b00100000;
            8'b10100011: signal <= 8'b00011110;
            8'b10100100: signal <= 8'b00011100;
            8'b10100101: signal <= 8'b00011010;
            8'b10100110: signal <= 8'b00011000;
            8'b10100111: signal <= 8'b00010111;
            8'b10101000: signal <= 8'b00010101;
            8'b10101001: signal <= 8'b00010011;
            8'b10101010: signal <= 8'b00010010;
            8'b10101011: signal <= 8'b00010000;
            8'b10101100: signal <= 8'b00001110;
            8'b10101101: signal <= 8'b00001101;
            8'b10101110: signal <= 8'b00001100;
            8'b10101111: signal <= 8'b00001010;
            8'b10110000: signal <= 8'b00001001;
            8'b10110001: signal <= 8'b00001000;
            8'b10110010: signal <= 8'b00000111;
            8'b10110011: signal <= 8'b00000110;
            8'b10110100: signal <= 8'b00000101;
            8'b10110101: signal <= 8'b00000100;
            8'b10110110: signal <= 8'b00000011;
            8'b10110111: signal <= 8'b00000011;
            8'b10111000: signal <= 8'b00000010;
            8'b10111001: signal <= 8'b00000001;
            8'b10111010: signal <= 8'b00000001;
            8'b10111011: signal <= 8'b00000000;
            8'b10111100: signal <= 8'b00000000;
            8'b10111101: signal <= 8'b00000000;
            8'b10111110: signal <= 8'b00000000;
            8'b10111111: signal <= 8'b00000000;
            8'b11000000: signal <= 8'b00000000;
            8'b11000001: signal <= 8'b00000000;
            8'b11000010: signal <= 8'b00000000;
            8'b11000011: signal <= 8'b00000000;
            8'b11000100: signal <= 8'b00000000;
            8'b11000101: signal <= 8'b00000000;
            8'b11000110: signal <= 8'b00000001;
            8'b11000111: signal <= 8'b00000001;
            8'b11001000: signal <= 8'b00000010;
            8'b11001001: signal <= 8'b00000011;
            8'b11001010: signal <= 8'b00000011;
            8'b11001011: signal <= 8'b00000100;
            8'b11001100: signal <= 8'b00000101;
            8'b11001101: signal <= 8'b00000110;
            8'b11001110: signal <= 8'b00000111;
            8'b11001111: signal <= 8'b00001000;
            8'b11010000: signal <= 8'b00001001;
            8'b11010001: signal <= 8'b00001010;
            8'b11010010: signal <= 8'b00001100;
            8'b11010011: signal <= 8'b00001101;
            8'b11010100: signal <= 8'b00001110;
            8'b11010101: signal <= 8'b00010000;
            8'b11010110: signal <= 8'b00010010;
            8'b11010111: signal <= 8'b00010011;
            8'b11011000: signal <= 8'b00010101;
            8'b11011001: signal <= 8'b00010111;
            8'b11011010: signal <= 8'b00011000;
            8'b11011011: signal <= 8'b00011010;
            8'b11011100: signal <= 8'b00011100;
            8'b11011101: signal <= 8'b00011110;
            8'b11011110: signal <= 8'b00100000;
            8'b11011111: signal <= 8'b00100011;
            8'b11100000: signal <= 8'b00100101;
            8'b11100001: signal <= 8'b00100111;
            8'b11100010: signal <= 8'b00101001;
            8'b11100011: signal <= 8'b00101100;
            8'b11100100: signal <= 8'b00101110;
            8'b11100101: signal <= 8'b00110000;
            8'b11100110: signal <= 8'b00110011;
            8'b11100111: signal <= 8'b00110101;
            8'b11101000: signal <= 8'b00111000;
            8'b11101001: signal <= 8'b00111011;
            8'b11101010: signal <= 8'b00111101;
            8'b11101011: signal <= 8'b01000000;
            8'b11101100: signal <= 8'b01000011;
            8'b11101101: signal <= 8'b01000101;
            8'b11101110: signal <= 8'b01001000;
            8'b11101111: signal <= 8'b01001011;
            8'b11110000: signal <= 8'b01001110;
            8'b11110001: signal <= 8'b01010001;
            8'b11110010: signal <= 8'b01010100;
            8'b11110011: signal <= 8'b01010111;
            8'b11110100: signal <= 8'b01011010;
            8'b11110101: signal <= 8'b01011101;
            8'b11110110: signal <= 8'b01100000;
            8'b11110111: signal <= 8'b01100011;
            8'b11111000: signal <= 8'b01100110;
            8'b11111001: signal <= 8'b01101001;
            8'b11111010: signal <= 8'b01101100;
            8'b11111011: signal <= 8'b01101111;
            8'b11111100: signal <= 8'b01110010;
            8'b11111101: signal <= 8'b01110101;
            8'b11111110: signal <= 8'b01111000;
            8'b11111111: signal <= 8'b01111011;
            default: signal <= 8'b00000000; // should never happen
        endcase
    end
endmodule
